module const_table#(

	parameter wordlength = 18,
	parameter LLR_wordlength = 19,
	parameter fraction = 10,
	parameter sym_num = 64,
	parameter bit_num = 6

)(
	input wire [2:0] 		Mode,
	output wire [wordlength-1:0] 	LUT_real_0, LUT_real_1, LUT_real_2, LUT_real_3, LUT_real_4, LUT_real_5, LUT_real_6, LUT_real_7, LUT_real_8, LUT_real_9, 
					LUT_real_10, LUT_real_11, LUT_real_12, LUT_real_13, LUT_real_14, LUT_real_15, LUT_real_16, LUT_real_17, LUT_real_18, LUT_real_19, 
					LUT_real_20, LUT_real_21, LUT_real_22, LUT_real_23, LUT_real_24, LUT_real_25, LUT_real_26, LUT_real_27, LUT_real_28, LUT_real_29, 
					LUT_real_30, LUT_real_31, LUT_real_32, LUT_real_33, LUT_real_34, LUT_real_35, LUT_real_36, LUT_real_37, LUT_real_38, LUT_real_39, 
					LUT_real_40, LUT_real_41, LUT_real_42, LUT_real_43, LUT_real_44, LUT_real_45, LUT_real_46, LUT_real_47, LUT_real_48, LUT_real_49, 
					LUT_real_50, LUT_real_51, LUT_real_52, LUT_real_53, LUT_real_54, LUT_real_55, LUT_real_56, LUT_real_57, LUT_real_58, LUT_real_59, 
					LUT_real_60, LUT_real_61, LUT_real_62, LUT_real_63,

	output wire [wordlength-1:0] 	LUT_imag_0, LUT_imag_1, LUT_imag_2, LUT_imag_3, LUT_imag_4, LUT_imag_5, LUT_imag_6, LUT_imag_7, LUT_imag_8, LUT_imag_9, 
					LUT_imag_10, LUT_imag_11, LUT_imag_12, LUT_imag_13, LUT_imag_14, LUT_imag_15, LUT_imag_16, LUT_imag_17, LUT_imag_18, LUT_imag_19, 
					LUT_imag_20, LUT_imag_21, LUT_imag_22, LUT_imag_23, LUT_imag_24, LUT_imag_25, LUT_imag_26, LUT_imag_27, LUT_imag_28, LUT_imag_29, 
					LUT_imag_30, LUT_imag_31, LUT_imag_32, LUT_imag_33, LUT_imag_34, LUT_imag_35, LUT_imag_36, LUT_imag_37, LUT_imag_38, LUT_imag_39, 
					LUT_imag_40, LUT_imag_41, LUT_imag_42, LUT_imag_43, LUT_imag_44, LUT_imag_45, LUT_imag_46, LUT_imag_47, LUT_imag_48, LUT_imag_49, 
					LUT_imag_50, LUT_imag_51, LUT_imag_52, LUT_imag_53, LUT_imag_54, LUT_imag_55, LUT_imag_56, LUT_imag_57, LUT_imag_58, LUT_imag_59, 
					LUT_imag_60, LUT_imag_61, LUT_imag_62, LUT_imag_63
);

assign LUT_real_0 = (Mode == 3'd1) ? 18'b000000001011010100 :
                      (Mode == 3'd2) ? 18'b000000001011010100 :
                      (Mode == 3'd3) ? 18'b000000001100110110 :
                      (Mode == 3'd4) ? 18'b111111110100100011 :
                      (Mode == 3'd5) ? 18'b000000001110110111 : 18'd0;

assign LUT_imag_0 = (Mode == 3'd1) ? 18'b000000001011010100 :
                      (Mode == 3'd2) ? 18'b000000001011010100 :
                      (Mode == 3'd3) ? 18'b000000001100110110 :
                      (Mode == 3'd4) ? 18'b000000010001001000 :
                      (Mode == 3'd5) ? 18'b000000001110110111 : 18'd0;

assign LUT_real_1 = (Mode == 3'd1) ? 18'b000000001011010100 :
                      (Mode == 3'd2) ? 18'b000000010000000000 :
                      (Mode == 3'd3) ? 18'b000000001100110110 :
                      (Mode == 3'd4) ? 18'b111111111011111110 :
                      (Mode == 3'd5) ? 18'b000000001110110111 : 18'd0;

assign LUT_imag_1 = (Mode == 3'd1) ? 18'b111111110100101011 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b111111110011001001 :
                      (Mode == 3'd4) ? 18'b000000010100001101 :
                      (Mode == 3'd5) ? 18'b111111110001001000 : 18'd0;

assign LUT_real_2 = (Mode == 3'd1) ? 18'b111111110100101011 :
                      (Mode == 3'd2) ? 18'b111111110000000000 :
                      (Mode == 3'd3) ? 18'b111111110011001001 :
                      (Mode == 3'd4) ? 18'b000000001011011100 :
                      (Mode == 3'd5) ? 18'b111111110001001000 : 18'd0;

assign LUT_imag_2 = (Mode == 3'd1) ? 18'b000000001011010100 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000001100110110 :
                      (Mode == 3'd4) ? 18'b000000010001001000 :
                      (Mode == 3'd5) ? 18'b000000001110110111 : 18'd0;

assign LUT_real_3 = (Mode == 3'd1) ? 18'b111111110100101011 :
                      (Mode == 3'd2) ? 18'b111111110100101011 :
                      (Mode == 3'd3) ? 18'b111111110011001001 :
                      (Mode == 3'd4) ? 18'b000000000100000001 :
                      (Mode == 3'd5) ? 18'b111111110001001000 : 18'd0;

assign LUT_imag_3 = (Mode == 3'd1) ? 18'b111111110100101011 :
                      (Mode == 3'd2) ? 18'b111111110100101011 :
                      (Mode == 3'd3) ? 18'b111111110011001001 :
                      (Mode == 3'd4) ? 18'b000000010100001101 :
                      (Mode == 3'd5) ? 18'b111111110001001000 : 18'd0;

assign LUT_real_4 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000010001100011 :
                      (Mode == 3'd4) ? 18'b111111111000100001 :
                      (Mode == 3'd5) ? 18'b000000000010010110 : 18'd0;

assign LUT_imag_4 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000010000000000 :
                      (Mode == 3'd3) ? 18'b000000000100101101 :
                      (Mode == 3'd4) ? 18'b000000000111011110 :
                      (Mode == 3'd5) ? 18'b000000010100111001 : 18'd0;

assign LUT_real_5 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000000001011010100 :
                      (Mode == 3'd3) ? 18'b000000010001100011 :
                      (Mode == 3'd4) ? 18'b111111111101010000 :
                      (Mode == 3'd5) ? 18'b000000000010010110 : 18'd0;

assign LUT_imag_5 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b111111110100101011 :
                      (Mode == 3'd3) ? 18'b111111111011010010 :
                      (Mode == 3'd4) ? 18'b000000001010001110 :
                      (Mode == 3'd5) ? 18'b111111101011000110 : 18'd0;

assign LUT_real_6 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b111111110100101011 :
                      (Mode == 3'd3) ? 18'b111111101110011100 :
                      (Mode == 3'd4) ? 18'b000000000111011110 :
                      (Mode == 3'd5) ? 18'b111111111101101001 : 18'd0;

assign LUT_imag_6 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000001011010100 :
                      (Mode == 3'd3) ? 18'b000000000100101101 :
                      (Mode == 3'd4) ? 18'b000000000111011110 :
                      (Mode == 3'd5) ? 18'b000000010100111001 : 18'd0;

assign LUT_real_7 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b111111101110011100 :
                      (Mode == 3'd4) ? 18'b000000000010101111 :
                      (Mode == 3'd5) ? 18'b111111111101101001 : 18'd0;

assign LUT_imag_7 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b111111110000000000 :
                      (Mode == 3'd3) ? 18'b111111111011010010 :
                      (Mode == 3'd4) ? 18'b000000001010001110 :
                      (Mode == 3'd5) ? 18'b111111101011000110 : 18'd0;

assign LUT_real_8 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000000000100101101 :
                      (Mode == 3'd4) ? 18'b111111101110110111 :
                      (Mode == 3'd5) ? 18'b000000010100111001 : 18'd0;

assign LUT_imag_8 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000010001100011 :
                      (Mode == 3'd4) ? 18'b000000001011011100 :
                      (Mode == 3'd5) ? 18'b000000000010010110 : 18'd0;

assign LUT_real_9 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000000000100101101 :
                      (Mode == 3'd4) ? 18'b111111101011110010 :
                      (Mode == 3'd5) ? 18'b000000010100111001 : 18'd0;

assign LUT_imag_9 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b111111101110011100 :
                      (Mode == 3'd4) ? 18'b000000000100000001 :
                      (Mode == 3'd5) ? 18'b111111111101101001 : 18'd0;

assign LUT_real_10 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b111111111011010010 :
                      (Mode == 3'd4) ? 18'b000000010001001000 :
                      (Mode == 3'd5) ? 18'b111111101011000110 : 18'd0;

assign LUT_imag_10 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000010001100011 :
                      (Mode == 3'd4) ? 18'b000000001011011100 :
                      (Mode == 3'd5) ? 18'b000000000010010110 : 18'd0;

assign LUT_real_11 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b111111111011010010 :
                      (Mode == 3'd4) ? 18'b000000010100001101 :
                      (Mode == 3'd5) ? 18'b111111101011000110 : 18'd0;

assign LUT_imag_11 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b111111101110011100 :
                      (Mode == 3'd4) ? 18'b000000000100000001 :
                      (Mode == 3'd5) ? 18'b111111111101101001 : 18'd0;

assign LUT_real_12 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000000000100000101 :
                      (Mode == 3'd4) ? 18'b111111110101110001 :
                      (Mode == 3'd5) ? 18'b000000000010000111 : 18'd0;

assign LUT_imag_12 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000100000101 :
                      (Mode == 3'd4) ? 18'b000000000010101111 :
                      (Mode == 3'd5) ? 18'b000000000010000111 : 18'd0;

assign LUT_real_13 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000000000100000101 :
                      (Mode == 3'd4) ? 18'b111111111101010111 :
                      (Mode == 3'd5) ? 18'b000000000010000111 : 18'd0;

assign LUT_imag_13 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b111111111011111010 :
                      (Mode == 3'd4) ? 18'b000000000010101000 :
                      (Mode == 3'd5) ? 18'b111111111101111000 : 18'd0;

assign LUT_real_14 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b111111111011111010 :
                      (Mode == 3'd4) ? 18'b000000001010001110 :
                      (Mode == 3'd5) ? 18'b111111111101111000 : 18'd0;

assign LUT_imag_14 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000100000101 :
                      (Mode == 3'd4) ? 18'b000000000010101111 :
                      (Mode == 3'd5) ? 18'b000000000010000111 : 18'd0;

assign LUT_real_15 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b111111111011111010 :
                      (Mode == 3'd4) ? 18'b000000000010101000 :
                      (Mode == 3'd5) ? 18'b111111111101111000 : 18'd0;

assign LUT_imag_15 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b111111111011111010 :
                      (Mode == 3'd4) ? 18'b000000000010101000 :
                      (Mode == 3'd5) ? 18'b111111111101111000 : 18'd0;

assign LUT_real_16 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111110100100011 :
                      (Mode == 3'd5) ? 18'b000000001011001100 : 18'd0;

assign LUT_imag_16 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111101110110111 :
                      (Mode == 3'd5) ? 18'b000000010001110011 : 18'd0;

assign LUT_real_17 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111111011111110 :
                      (Mode == 3'd5) ? 18'b000000001011001100 : 18'd0;

assign LUT_imag_17 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111101011110010 :
                      (Mode == 3'd5) ? 18'b111111101110001100 : 18'd0;

assign LUT_real_18 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000001011011100 :
                      (Mode == 3'd5) ? 18'b111111110100110011 : 18'd0;

assign LUT_imag_18 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111101110110111 :
                      (Mode == 3'd5) ? 18'b000000010001110011 : 18'd0;

assign LUT_real_19 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000000100000001 :
                      (Mode == 3'd5) ? 18'b111111110100110011 : 18'd0;

assign LUT_imag_19 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111101011110010 :
                      (Mode == 3'd5) ? 18'b111111101110001100 : 18'd0;

assign LUT_real_20 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111111000100001 :
                      (Mode == 3'd5) ? 18'b000000000110111100 : 18'd0;

assign LUT_imag_20 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111000100001 :
                      (Mode == 3'd5) ? 18'b000000010011110110 : 18'd0;

assign LUT_real_21 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111111101010000 :
                      (Mode == 3'd5) ? 18'b000000000110111100 : 18'd0;

assign LUT_imag_21 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111110101110001 :
                      (Mode == 3'd5) ? 18'b111111101100001001 : 18'd0;

assign LUT_real_22 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000000111011110 :
                      (Mode == 3'd5) ? 18'b111111111001000011 : 18'd0;

assign LUT_imag_22 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111000100001 :
                      (Mode == 3'd5) ? 18'b000000010011110110 : 18'd0;

assign LUT_real_23 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000000010101111 :
                      (Mode == 3'd5) ? 18'b111111111001000011 : 18'd0;

assign LUT_imag_23 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111110101110001 :
                      (Mode == 3'd5) ? 18'b111111101100001001 : 18'd0;

assign LUT_real_24 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111101110110111 :
                      (Mode == 3'd5) ? 18'b000000001100110000 : 18'd0;

assign LUT_imag_24 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111110100100011 :
                      (Mode == 3'd5) ? 18'b000000000010000001 : 18'd0;

assign LUT_real_25 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111101011110010 :
                      (Mode == 3'd5) ? 18'b000000001100110000 : 18'd0;

assign LUT_imag_25 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111011111110 :
                      (Mode == 3'd5) ? 18'b111111111101111110 : 18'd0;

assign LUT_real_26 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000010001001000 :
                      (Mode == 3'd5) ? 18'b111111110011001111 : 18'd0;

assign LUT_imag_26 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111110100100011 :
                      (Mode == 3'd5) ? 18'b000000000010000001 : 18'd0;

assign LUT_real_27 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000010100001101 :
                      (Mode == 3'd5) ? 18'b111111110011001111 : 18'd0;

assign LUT_imag_27 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111011111110 :
                      (Mode == 3'd5) ? 18'b111111111101111110 : 18'd0;

assign LUT_real_28 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111110101110001 :
                      (Mode == 3'd5) ? 18'b000000000110111101 : 18'd0;

assign LUT_imag_28 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111101010000 :
                      (Mode == 3'd5) ? 18'b000000000001110111 : 18'd0;

assign LUT_real_29 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b111111111101010111 :
                      (Mode == 3'd5) ? 18'b000000000110111101 : 18'd0;

assign LUT_imag_29 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111101010111 :
                      (Mode == 3'd5) ? 18'b111111111110001000 : 18'd0;

assign LUT_real_30 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000001010001110 :
                      (Mode == 3'd5) ? 18'b111111111001000010 : 18'd0;

assign LUT_imag_30 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111101010000 :
                      (Mode == 3'd5) ? 18'b000000000001110111 : 18'd0;

assign LUT_real_31 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000000000010101000 :
                      (Mode == 3'd5) ? 18'b111111111001000010 : 18'd0;

assign LUT_imag_31 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b111111111101010111 :
                      (Mode == 3'd5) ? 18'b111111111110001000 : 18'd0;

assign LUT_real_32 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000010001110011 : 18'd0;

assign LUT_imag_32 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001011001100 : 18'd0;

assign LUT_real_33 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000010001110011 : 18'd0;

assign LUT_imag_33 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110100110011 : 18'd0;

assign LUT_real_34 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111101110001100 : 18'd0;

assign LUT_imag_34 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001011001100 : 18'd0;

assign LUT_real_35 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111101110001100 : 18'd0;

assign LUT_imag_35 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110100110011 : 18'd0;

assign LUT_real_36 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000010000001 : 18'd0;

assign LUT_imag_36 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001100110000 : 18'd0;

assign LUT_real_37 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000010000001 : 18'd0;

assign LUT_imag_37 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110011001111 : 18'd0;

assign LUT_real_38 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111101111110 : 18'd0;

assign LUT_imag_38 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001100110000 : 18'd0;

assign LUT_real_39 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111101111110 : 18'd0;

assign LUT_imag_39 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110011001111 : 18'd0;

assign LUT_real_40 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000010011110110 : 18'd0;

assign LUT_imag_40 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000110111100 : 18'd0;

assign LUT_real_41 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000010011110110 : 18'd0;

assign LUT_imag_41 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111001000011 : 18'd0;

assign LUT_real_42 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111101100001001 : 18'd0;

assign LUT_imag_42 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000110111100 : 18'd0;

assign LUT_real_43 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111101100001001 : 18'd0;

assign LUT_imag_43 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111001000011 : 18'd0;

assign LUT_real_44 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000001110111 : 18'd0;

assign LUT_imag_44 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000110111101 : 18'd0;

assign LUT_real_45 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000001110111 : 18'd0;

assign LUT_imag_45 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111001000010 : 18'd0;

assign LUT_real_46 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111110001000 : 18'd0;

assign LUT_imag_46 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000110111101 : 18'd0;

assign LUT_real_47 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111110001000 : 18'd0;

assign LUT_imag_47 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111001000010 : 18'd0;

assign LUT_real_48 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000001001001000 : 18'd0;

assign LUT_imag_48 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001001001000 : 18'd0;

assign LUT_real_49 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000001001001000 : 18'd0;

assign LUT_imag_49 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110110110111 : 18'd0;

assign LUT_real_50 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111110110110111 : 18'd0;

assign LUT_imag_50 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001001001000 : 18'd0;

assign LUT_real_51 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111110110110111 : 18'd0;

assign LUT_imag_51 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110110110111 : 18'd0;

assign LUT_real_52 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000101110111 : 18'd0;

assign LUT_imag_52 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001011100000 : 18'd0;

assign LUT_real_53 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000101110111 : 18'd0;

assign LUT_imag_53 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110100011111 : 18'd0;

assign LUT_real_54 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111010001000 : 18'd0;

assign LUT_imag_54 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000001011100000 : 18'd0;

assign LUT_real_55 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111010001000 : 18'd0;

assign LUT_imag_55 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111110100011111 : 18'd0;

assign LUT_real_56 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000001011100000 : 18'd0;

assign LUT_imag_56 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000101110111 : 18'd0;

assign LUT_real_57 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000001011100000 : 18'd0;

assign LUT_imag_57 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111010001000 : 18'd0;

assign LUT_real_58 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111110100011111 : 18'd0;

assign LUT_imag_58 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000101110111 : 18'd0;

assign LUT_real_59 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111110100011111 : 18'd0;

assign LUT_imag_59 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111010001000 : 18'd0;

assign LUT_real_60 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000101000110 : 18'd0;

assign LUT_imag_60 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000101000110 : 18'd0;

assign LUT_real_61 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b000000000101000110 : 18'd0;

assign LUT_imag_61 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111010111001 : 18'd0;

assign LUT_real_62 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111010111001 : 18'd0;

assign LUT_imag_62 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b000000000101000110 : 18'd0;

assign LUT_real_63 = (Mode == 3'd1) ? 18'b000001100000000000 :
                      (Mode == 3'd2) ? 18'b000001010000000000 :
                      (Mode == 3'd3) ? 18'b000001010000000000 :
                      (Mode == 3'd4) ? 18'b000001010000000000 :
                      (Mode == 3'd5) ? 18'b111111111010111001 : 18'd0;

assign LUT_imag_63 = (Mode == 3'd1) ? 18'b000000000000000000 :
                      (Mode == 3'd2) ? 18'b000000000000000000 :
                      (Mode == 3'd3) ? 18'b000000000000000000 :
                      (Mode == 3'd4) ? 18'b000000000000000000 :
                      (Mode == 3'd5) ? 18'b111111111010111001 : 18'd0;
	      
endmodule
