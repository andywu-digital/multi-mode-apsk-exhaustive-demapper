`define WORDLENGTH 18 //Q8.10
module Vectoring_Mode(clk, rst_n, en, x_i, y_i, valid, z_o);

input   clk, rst_n, en;
input   signed  [`WORDLENGTH-1:0] x_i, y_i;

output  reg valid;
output  reg signed  [`WORDLENGTH-1:0] z_o;

// ===================== //
// Prerotation 
// ===================== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]    xi_inv, yi_inv, x_pre, y_pre, z_pre, x_pre_o, y_pre_o, z_pre_o;
wire    angle_pre, pre_rot;   
// -------------- //
assign {angle_pre, pre_rot} = {y_i[`WORDLENGTH-1], x_i[`WORDLENGTH-1]}; 

assign xi_inv = -x_i;
assign yi_inv = -y_i;

assign x_pre = (angle_pre)? yi_inv:y_i;
assign y_pre = (angle_pre)? x_i:xi_inv;
assign z_pre = (angle_pre)? 18'h3f9b7:18'h00648; //pi/2

assign x_pre_o = (pre_rot)? x_pre:x_i;
assign y_pre_o = (pre_rot)? y_pre:y_i;
assign z_pre_o = (pre_rot)? z_pre:{`WORDLENGTH{1'd0}};

// ========== //
// Stage 0
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   x_s0_inv, y_s0_inv, x_s0_sel, y_s0_sel, z_s0_sel, x_s0_o, y_s0_o, z_s0_o;
wire    angle_0;
// -------------- //
assign angle_0 = y_pre_o[`WORDLENGTH-1];

assign x_s0_inv = -x_pre_o;
assign y_s0_inv = -y_pre_o;

assign x_s0_sel = (angle_0)? y_s0_inv:y_pre_o;
assign y_s0_sel = (angle_0)? x_pre_o:x_s0_inv;
assign z_s0_sel = (angle_0)? 18'h3fcdc:18'h00324; //atan(2^(-0))

assign x_s0_o = x_pre_o + x_s0_sel;
assign y_s0_o = y_pre_o + y_s0_sel;
assign z_s0_o = z_pre_o + z_s0_sel;

// ========== //
// Stage 1
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   x_s1_inv, y_s1_inv, x_s1_sel, y_s1_sel, z_s1_sel, x_s1_shf, y_s1_shf;
wire    signed  [`WORDLENGTH-1:0]   x_s1_o, y_s1_o, z_s1_o;
wire    angle_1;
// -------------- //
assign angle_1 = y_s0_o[`WORDLENGTH-1];

assign x_s1_inv = -x_s0_o;
assign y_s1_inv = -y_s0_o;

assign x_s1_sel = (angle_1)? y_s1_inv:y_s0_o;
assign y_s1_sel = (angle_1)? x_s0_o:x_s1_inv;
assign z_s1_sel = (angle_1)? 18'h3fe26:18'h001da; //atan(2^(-1))

assign x_s1_shf = x_s1_sel>>>1;
assign y_s1_shf = y_s1_sel>>>1;

assign x_s1_o = x_s0_o + x_s1_shf;
assign y_s1_o = y_s0_o + y_s1_shf;
assign z_s1_o = z_s0_o + z_s1_sel;

// ========== //
// Stage 2
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   x_s2_inv, y_s2_inv, x_s2_sel, y_s2_sel, z_s2_sel, x_s2_shf, y_s2_shf;
wire    signed  [`WORDLENGTH-1:0]   x_s2_o, y_s2_o, z_s2_o;
wire    angle_2;
// -------------- //
assign angle_2 = y_s1_o[`WORDLENGTH-1];

assign x_s2_inv = -x_s1_o;
assign y_s2_inv = -y_s1_o;

assign x_s2_sel = (angle_2)? y_s2_inv:y_s1_o;
assign y_s2_sel = (angle_2)? x_s1_o:x_s2_inv;
assign z_s2_sel = (angle_2)? 18'h3ff06:18'h000fa; //atan(2^(-2))

assign x_s2_shf = x_s2_sel>>>2;
assign y_s2_shf = y_s2_sel>>>2;

assign x_s2_o = x_s1_o + x_s2_shf;
assign y_s2_o = y_s1_o + y_s2_shf;
assign z_s2_o = z_s1_o + z_s2_sel;

// ========== //
// Stage 3
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   x_s3_inv, y_s3_inv, x_s3_sel, y_s3_sel, z_s3_sel, x_s3_shf, y_s3_shf;
wire    signed  [`WORDLENGTH-1:0]   x_s3_o, y_s3_o, z_s3_o;
wire    angle_3;
// -------------- //
assign angle_3 = y_s2_o[`WORDLENGTH-1];

assign x_s3_inv = -x_s2_o;
assign y_s3_inv = -y_s2_o;

assign x_s3_sel = (angle_3)? y_s3_inv:y_s2_o;
assign y_s3_sel = (angle_3)? x_s2_o:x_s3_inv;
assign z_s3_sel = (angle_3)? 18'h3ff81:18'h0007f; //atan(2^(-3))

assign x_s3_shf = x_s3_sel>>>3;
assign y_s3_shf = y_s3_sel>>>3;

assign x_s3_o = x_s2_o + x_s3_shf;
assign y_s3_o = y_s2_o + y_s3_shf;
assign z_s3_o = z_s2_o + z_s3_sel;

// ========== //
// Stage 4
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   x_s4_inv, y_s4_inv, x_s4_sel, y_s4_sel, z_s4_sel, x_s4_shf, y_s4_shf;
wire    signed  [`WORDLENGTH-1:0]   x_s4_o, y_s4_o, z_s4_o;
wire    angle_4;
// -------------- //
assign angle_4 = y_s3_o[`WORDLENGTH-1];

assign x_s4_inv = -x_s3_o;
assign y_s4_inv = -y_s3_o;

assign x_s4_sel = (angle_4)? y_s4_inv:y_s3_o;
assign y_s4_sel = (angle_4)? x_s3_o:x_s4_inv;
assign z_s4_sel = (angle_4)? 18'h3ffc1:18'h0003f; //atan(2^(-4))

assign x_s4_shf = x_s4_sel>>>4;
assign y_s4_shf = y_s4_sel>>>4;

assign x_s4_o = x_s3_o + x_s4_shf;
assign y_s4_o = y_s3_o + y_s4_shf;
assign z_s4_o = z_s3_o + z_s4_sel;

// ========== //
// Stage 5
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   x_s5_inv, y_s5_sel, z_s5_sel, y_s5_shf;
wire    signed  [`WORDLENGTH-1:0]    y_s5_o, z_s5_o;
wire    angle_5;
// -------------- //
assign angle_5 = y_s4_o[`WORDLENGTH-1];

assign x_s5_inv = -x_s4_o;



assign y_s5_sel = (angle_5)? x_s4_o:x_s5_inv;
assign z_s5_sel = (angle_5)? 18'h3ffe1:18'h0001f; //atan(2^(-5))


assign y_s5_shf = y_s5_sel>>>5;


assign y_s5_o = y_s4_o + y_s5_shf;
assign z_s5_o = z_s4_o + z_s5_sel;

// ========== //
// Stage 6
// ========== //
// --- Signal --- //
wire    signed  [`WORDLENGTH-1:0]   z_s6_sel;
wire    signed  [`WORDLENGTH-1:0]   z_s6_o;
wire    angle_6;
// -------------- //
assign angle_6 = y_s5_o[`WORDLENGTH-1];

assign z_s6_sel = (angle_6)? 18'b111111111111110001:18'b000000000000001111; //atan(2^(-6))

assign z_s6_o = z_s5_o + z_s6_sel;

// ========== //
// Output
// ========== //
always@(posedge clk or negedge rst_n)
    if(!rst_n) 
        valid <= 1'b0;
    else
        valid <= en;

always@(posedge clk or negedge rst_n)
    if(!rst_n) 
        z_o <= {`WORDLENGTH{1'd0}};
    else 
        z_o <= z_s6_o;

endmodule
